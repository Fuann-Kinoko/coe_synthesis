`define regwrite_ON 		1'b1
`define regwrite_OFF        1'b0

`define regdst_RD           1'b1
`define regdst_RT           1'b0

`define alusrc_IMM          1'b1
`define alusrc_RD           1'b0

`define branch_ON           1'b1
`define branch_OFF          1'b0

`define bal_ON              1'b1
`define bal_OFF             1'b0

`define memWrite_ON         1'b1
`define memWrite_OFF        1'b0

`define memToReg_MEM        1'b1
`define memToReg_ALU        1'b0

`define jump_ON             1'b1
`define jump_OFF            1'b0

`define jal_ON              1'b1
`define jal_OFF             1'b0